module evenparity(a,z);//?????
input[7:0] a;//8?? a
output[8:0] z;//9?? z
reg [8:0] z;//9?? ???? z
integer n,i;//n:1? ?? ???
always@(a)//a? ????
begin
n=0;//n? ???
for(i=0;i<8;i=i+1)begin
 z[i+1]=a[i];//z[1~8]=a[0~7]
if(a[i]==1) n=n+1;//n???
end
if(n%2==1) z[0]=1;//??
else  z[0]=0;//??
end
endmodule
