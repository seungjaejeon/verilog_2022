
module clock(t);
output t;

reg t;

endmodule