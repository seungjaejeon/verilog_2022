module alarm_clk(Clock_1Sec, Reset, LoadTime, LoadAlm,
AlarmEnable, Set_AM_PM, Alarm_AM_PM_In,
SetSecs, SetMins, AlarmMinsIn, SetHours, AlarmHoursIn,
AM_PM, Alarm, Secs_C, Mins_C, Hours_C);
input Clock_1Sec, Reset, LoadTime, LoadAlm, Set_AM_PM,
Alarm_AM_PM_In,AlarmEnable;
input[5:0] SetSecs, SetMins,AlarmMinsIn;
input[3:0] SetHours, AlarmHoursIn;
output AM_PM, Alarm;
output[5:0] Secs_C, Mins_C;
output[3:0] Hours_C;
reg AM_PM, Alarm,Alarm_AM_PM;
reg[5:0] Secs_C, Mins_C, AlarmMin;
reg[3:0] Hours_C,AlarmHour;

always@(negedge Reset)//???
begin
if(!Reset)//Reset? 0??
begin
AM_PM<=0;
Secs_C<=0;
Mins_C<=0;
Hours_C<=12;
AlarmMin<=0;
AlarmHour<=0;
Alarm_AM_PM<=0;
Alarm<=0;
end
end
always@(posedge Clock_1Sec)
begin
if(Reset)
begin
if(LoadTime==1)//?? ???(LoadTime? 1??)
begin//?? ? ??
	AM_PM<=Set_AM_PM;
	Secs_C<=SetSecs;
	Mins_C<=SetMins;
	Hours_C<=SetHours;
end
else//LoadTime? 0??
begin
Secs_C<=Secs_C+1;//1? ??
	if(Secs_C==59)//Secs_C=59?? 
	begin
	Secs_C<=0;//Secs_C? 0?? ??
	Mins_C<=Mins_C+1;//Mins_C? 1 ??
		if(Mins_C==59)//Mins_C? 59??
		begin
		Mins_C<=0;//Mins_C? 0?? ??
		Hours_C<=Hours_C+1;//Hours_C? 1??
			if(Hours_C==11) AM_PM<=~AM_PM;//Hours_C? 11?? ??????(11? 59? 59??? ??)
		else if(Hours_C==12) Hours_C<=1;//Hours_C? 12?? 1? ??
		end
	end
end
if(LoadAlm)//?? ??(LoadAlm? 1??)
	begin//???? ??? ???? ??
	AlarmMin<=AlarmMinsIn;
	AlarmHour<=AlarmHoursIn;
	Alarm_AM_PM<=Alarm_AM_PM_In;
	end
else//LoadAlm? 0??
begin
if(AlarmEnable)//ALarmEnable=1?? (??? ?? ? ??)
begin
	if(AlarmMin==0)//????? ?? 0? ?
	begin
		if(AlarmHour==12)//????? ?? 12??
		begin//AlarmHour=12,AlarmMin=0??
//??? ????? ?? ????? ??? ???? ????? 1?? ?? 59? ?? 59??? Alarm=1??
			if(AM_PM!=Alarm_AM_PM && Hours_C==AlarmHour-1 &&
			Mins_C==59 && Secs_C==59) Alarm<=1;
		end
		else if(AlarmHour==1)//????? 1? 00?? ??????
		begin
		if(AM_PM==Alarm_AM_PM && Hours_C==12 &&
		Mins_C==59 && Secs_C==59) Alarm<=1;
		end
		else//AlarmHour=12? ??? AlarmMin=0?? 
//??? ????? ?? ????? ?? ???? ????? 1?? ?? 59? ?? 59??? ALarm=1??
		if(AM_PM==Alarm_AM_PM && Hours_C==AlarmHour-1 &&
		Mins_C==59 && Secs_C==59) Alarm<=1;
	end
//AlarmHour=12, AlarmMin=0? ??? ??? ????? ?? ????? ?? ???? ???? ?? ?? 1???? ?? 59??? ALarm=1??
	else if(AM_PM==Alarm_AM_PM && Hours_C==AlarmHour
	&& Mins_C==AlarmMin-1 && Secs_C==59) Alarm<=1; 
end
if(Alarm==1)//Alarm=1??
begin//Secs_C? 59?? ?? Alarm? 0? ????? ? 1?? ???? ??.
if(Secs_C==59) Alarm<=0;
end
end
end
end
endmodule